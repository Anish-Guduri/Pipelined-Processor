module ALU_Stage(



);
endmodule