module ALU_Stage(
    input [9:0] input_EX_PC,
    input [31:0] EX_branchTarget,
    input [31:0] Operand_EX_A,
    input [31:0] Operand_EX_B,
    input [31:0] Operand_EX_2,
    input [31:0] input_EX_IR,
    output reg[31:0] output_EX_PC,
    output reg[31:0] ALU_Result,
    output reg[31:0] op2,
    output reg[31:0] output_EX_IR

);

always @(*) begin

        
end

endmodule